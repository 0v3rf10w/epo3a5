configuration buf_5_behaviour_cfg of buf_5 is
   for behaviour
   end for;
end buf_5_behaviour_cfg;


