configuration reg_4_behaviour_cfg of reg_4 is
   for behaviour
   end for;
end reg_4_behaviour_cfg;


