configuration spi_structural_cfg of spi is
   for structural
   end for;
end spi_structural_cfg;


