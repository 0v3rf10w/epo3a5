configuration klokdeler_behavioural_cfg of klokdeler is
   for behavioural
      for all: dff use configuration work.dff_behavioural_cfg;
      end for;
   end for;
end klokdeler_behavioural_cfg;


