configuration spi_slave_extracted_cfg of spi_slave is
   for extracted
   end for;
end spi_slave_extracted_cfg;


