configuration shift_reg_behaviour_cfg of shift_reg is
   for behaviour
   end for;
end shift_reg_behaviour_cfg;


