<<<<<<< HEAD
library IEEE;
use IEEE.std_logic_1164.ALL;

entity stream is
   port(IN_0 :in    std_logic;
        IN_1 :in    std_logic;
        OUT_0:out   std_logic;
        OUT_1:out   std_logic;
        E    :in    std_logic);
=======
library IEEE;
use IEEE.std_logic_1164.ALL;

entity stream is
   port(IN_0 :in    std_logic;
        IN_1 :in    std_logic;
        OUT_0:out   std_logic;
        OUT_1:out   std_logic;
        E    :in    std_logic);
>>>>>>> origin/master
end stream;


