configuration reg_5_behaviour_cfg of reg_5 is
   for behaviour
   end for;
end reg_5_behaviour_cfg;


