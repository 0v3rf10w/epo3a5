configuration buf_9_behaviour_cfg of buf_9 is
   for behaviour
   end for;
end buf_9_behaviour_cfg;


