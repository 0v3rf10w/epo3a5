configuration rom_behavioural_cfg of rom is
   for behavioural
   end for;
end rom_behavioural_cfg;


