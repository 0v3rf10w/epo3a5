configuration buf_6_behaviour_cfg of buf_6 is
   for behaviour
   end for;
end buf_6_behaviour_cfg;


