library IEEE;
use IEEE.std_logic_1164.ALL;

entity tbuf_tb is
end tbuf_tb;


