configuration counter_synthesised_cfg of counter is
   for synthesised
   end for;
end counter_synthesised_cfg;


