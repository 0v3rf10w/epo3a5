library IEEE;
use IEEE.std_logic_1164.ALL;

entity deler is
   port(clk      :in    std_logic;
        deler_out:out   std_logic);
end deler;


