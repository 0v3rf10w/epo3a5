configuration buf_7_behaviour_cfg of buf_7 is
   for behaviour
   end for;
end buf_7_behaviour_cfg;


