library IEEE;
use IEEE.std_logic_1164.ALL;

entity blackbox_tb is
end blackbox_tb;


