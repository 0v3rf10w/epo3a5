configuration reg_9_behaviour_cfg of reg_9 is
   for behaviour
   end for;
end reg_9_behaviour_cfg;


