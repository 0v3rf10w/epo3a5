configuration tb_behavioral_cfg of tb is
   for behavioral
      for all: calculator use configuration work.calculator_behaviour_cfg;
      end for;
   end for;
end tb_behavioral_cfg;


