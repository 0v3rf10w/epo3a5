configuration decoder_behaviour_cfg of decoder is
   for behaviour
   end for;
end decoder_behaviour_cfg;


