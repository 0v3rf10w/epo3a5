configuration buf_3_behaviour_cfg of buf_3 is
   for behaviour
   end for;
end buf_3_behaviour_cfg;


