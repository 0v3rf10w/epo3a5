configuration tb_behavioural_synt_cfg of tb is
   for behavioural
      for all: klokdeler use configuration work.klokdeler_behavioural_cfg;
      end for;
   end for;
end tb_behavioural_synt_cfg;


