configuration control_synthesised_cfg of control is
   for synthesised
   end for;
end control_synthesised_cfg;


