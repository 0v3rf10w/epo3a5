configuration shift_reg_synthesised_cfg of shift_reg is
   for synthesised
   end for;
end shift_reg_synthesised_cfg;


