library IEEE;
use IEEE.std_logic_1164.ALL;

entity iv is
   port(A:in    std_logic;
        Y:out    std_logic);
end iv;


