
library ieee,CellsLib;

use ieee.std_logic_1164.all;
use CellsLib.CellsLib_DECL_PACK.all;

architecture synthesised of rom is

   component iv110
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   component no210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component na210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component na310
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component no310
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   signal n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820 : std_logic;

begin
   
   U429 : na310 port map( A => n417, B => n418, C => n419, Y => rom_d(9));
   U430 : no310 port map( A => n420, B => n421, C => n422, Y => n419);
   U431 : no210 port map( A => n423, B => n424, Y => n420);
   U432 : no210 port map( A => n425, B => n426, Y => n423);
   U433 : no210 port map( A => n427, B => n428, Y => n417);
   U434 : na310 port map( A => n429, B => n430, C => n431, Y => rom_d(8));
   U435 : iv110 port map( A => n432, Y => n431);
   U436 : na210 port map( A => n433, B => n434, Y => n432);
   U437 : no310 port map( A => n435, B => n436, C => n437, Y => n434);
   U438 : no310 port map( A => n438, B => n439, C => n440, Y => n433);
   U439 : no310 port map( A => n441, B => n422, C => n442, Y => n430);
   U440 : no210 port map( A => n443, B => n444, Y => n442);
   U441 : no210 port map( A => n445, B => n446, Y => n443);
   U442 : na210 port map( A => n447, B => n448, Y => n441);
   U443 : na210 port map( A => n449, B => n450, Y => n448);
   U444 : na210 port map( A => n451, B => n452, Y => n447);
   U445 : no310 port map( A => n453, B => n454, C => n455, Y => n429);
   U446 : no210 port map( A => n456, B => n457, Y => n455);
   U447 : no210 port map( A => n458, B => n459, Y => n454);
   U448 : na310 port map( A => n460, B => n461, C => n462, Y => rom_d(7));
   U449 : no310 port map( A => n463, B => n464, C => n465, Y => n462);
   U450 : no210 port map( A => n466, B => n424, Y => n465);
   U451 : no210 port map( A => n467, B => n468, Y => n464);
   U452 : no210 port map( A => n469, B => n470, Y => n467);
   U453 : na210 port map( A => n471, B => n472, Y => n461);
   U454 : iv110 port map( A => n473, Y => n460);
   U455 : na210 port map( A => n474, B => n475, Y => rom_d(6));
   U456 : no310 port map( A => n476, B => n422, C => n477, Y => n475);
   U457 : no210 port map( A => n478, B => n479, Y => n477);
   U458 : no210 port map( A => n480, B => n481, Y => n478);
   U459 : no210 port map( A => n482, B => n466, Y => n422);
   U460 : no210 port map( A => n483, B => n424, Y => n476);
   U461 : no310 port map( A => n484, B => n485, C => n486, Y => n474);
   U462 : no210 port map( A => n466, B => n487, Y => n486);
   U463 : no210 port map( A => n488, B => n459, Y => n485);
   U464 : na310 port map( A => n489, B => n490, C => n491, Y => rom_d(5));
   U465 : no310 port map( A => n492, B => n493, C => n494, Y => n491);
   U466 : no210 port map( A => n487, B => n495, Y => n494);
   U467 : no210 port map( A => n456, B => n466, Y => n492);
   U468 : no210 port map( A => n496, B => n427, Y => n489);
   U469 : na310 port map( A => n497, B => n498, C => n499, Y => n427);
   U470 : no310 port map( A => n473, B => n500, C => n501, Y => n499);
   U471 : na310 port map( A => n502, B => n503, C => n504, Y => n473);
   U472 : no210 port map( A => n505, B => n506, Y => n504);
   U473 : no210 port map( A => n507, B => n508, Y => n506);
   U474 : na210 port map( A => n509, B => n510, Y => n503);
   U475 : na210 port map( A => n450, B => n511, Y => n498);
   U476 : no210 port map( A => n512, B => n513, Y => n497);
   U477 : iv110 port map( A => n514, Y => n513);
   U478 : na210 port map( A => n426, B => n480, Y => n514);
   U479 : na210 port map( A => n515, B => n459, Y => n426);
   U480 : no210 port map( A => n516, B => n456, Y => n512);
   U481 : iv110 port map( A => n517, Y => n516);
   U482 : na310 port map( A => n518, B => n519, C => n520, Y => rom_d(4));
   U483 : no310 port map( A => n521, B => n522, C => n523, Y => n520);
   U484 : no210 port map( A => n466, B => n468, Y => n523);
   U485 : no210 port map( A => n524, B => n457, Y => n522);
   U486 : iv110 port map( A => n525, Y => n521);
   U487 : no210 port map( A => n526, B => n421, Y => n525);
   U488 : no210 port map( A => n482, B => n527, Y => n526);
   U489 : iv110 port map( A => n528, Y => n519);
   U490 : no210 port map( A => n484, B => n529, Y => n518);
   U491 : na310 port map( A => n530, B => n531, C => n532, Y => n484);
   U492 : no310 port map( A => n533, B => n493, C => n505, Y => n532);
   U493 : no210 port map( A => n534, B => n507, Y => n533);
   U494 : na210 port map( A => n535, B => n536, Y => n531);
   U495 : iv110 port map( A => n537, Y => n530);
   U496 : na310 port map( A => n538, B => n539, C => n540, Y => rom_d(3));
   U497 : no310 port map( A => n541, B => n542, C => n543, Y => n540);
   U498 : no210 port map( A => n457, B => n507, Y => n542);
   U499 : na210 port map( A => n544, B => n545, Y => n541);
   U500 : na210 port map( A => n510, B => n546, Y => n545);
   U501 : na210 port map( A => n515, B => n466, Y => n546);
   U502 : no210 port map( A => n436, B => n537, Y => n539);
   U503 : na310 port map( A => n547, B => n548, C => n549, Y => n436);
   U504 : no310 port map( A => n550, B => n551, C => n552, Y => n549);
   U505 : no210 port map( A => n553, B => n534, Y => n551);
   U506 : na210 port map( A => n452, B => n446, Y => n548);
   U507 : iv110 port map( A => n554, Y => n446);
   U508 : no210 port map( A => n555, B => n556, Y => n547);
   U509 : no210 port map( A => n557, B => n558, Y => n556);
   U510 : no210 port map( A => n559, B => n509, Y => n557);
   U511 : no210 port map( A => n560, B => n561, Y => n555);
   U512 : no210 port map( A => n469, B => n562, Y => n560);
   U513 : no210 port map( A => n563, B => n564, Y => n538);
   U514 : na310 port map( A => n565, B => n566, C => n567, Y => rom_d(2));
   U515 : no310 port map( A => n568, B => n569, C => n570, Y => n567);
   U516 : no210 port map( A => n571, B => n507, Y => n570);
   U517 : no210 port map( A => n424, B => n508, Y => n569);
   U518 : iv110 port map( A => n572, Y => n568);
   U519 : no310 port map( A => n573, B => n574, C => n575, Y => n572);
   U520 : no210 port map( A => n561, B => n576, Y => n575);
   U521 : no210 port map( A => n558, B => n577, Y => n574);
   U522 : no210 port map( A => n468, B => n578, Y => n573);
   U523 : no310 port map( A => n550, B => n579, C => n580, Y => n566);
   U524 : no210 port map( A => n581, B => n457, Y => n579);
   U525 : na310 port map( A => n582, B => n583, C => n584, Y => n550);
   U526 : no210 port map( A => n493, B => n421, Y => n584);
   U527 : no210 port map( A => n456, B => n585, Y => n421);
   U528 : na210 port map( A => n469, B => n586, Y => n583);
   U529 : na210 port map( A => n559, B => n536, Y => n582);
   U530 : no210 port map( A => n440, B => n563, Y => n565);
   U531 : iv110 port map( A => n587, Y => n563);
   U532 : na310 port map( A => n588, B => n589, C => n590, Y => n440);
   U533 : iv110 port map( A => n591, Y => n590);
   U534 : na210 port map( A => n449, B => n592, Y => n589);
   U535 : na310 port map( A => n593, B => n594, C => n595, Y => rom_d(1));
   U536 : iv110 port map( A => n596, Y => n595);
   U537 : na310 port map( A => n597, B => n490, C => n587, Y => n596);
   U538 : no210 port map( A => n598, B => n599, Y => n587);
   U539 : no310 port map( A => n600, B => n601, C => n435, Y => n597);
   U540 : na210 port map( A => n602, B => n603, Y => n435);
   U541 : no310 port map( A => n604, B => n605, C => n606, Y => n603);
   U542 : no210 port map( A => n607, B => n558, Y => n606);
   U543 : no210 port map( A => n608, B => n515, Y => n605);
   U544 : no210 port map( A => n536, B => n609, Y => n608);
   U545 : na210 port map( A => n610, B => n611, Y => n604);
   U546 : na210 port map( A => n449, B => n612, Y => n611);
   U547 : na210 port map( A => n469, B => n471, Y => n610);
   U548 : no310 port map( A => n613, B => n614, C => n580, Y => n602);
   U549 : na310 port map( A => n615, B => n616, C => n617, Y => n580);
   U550 : no210 port map( A => n618, B => n619, Y => n617);
   U551 : no210 port map( A => n620, B => n558, Y => n619);
   U552 : no210 port map( A => n621, B => n561, Y => n618);
   U553 : no210 port map( A => n622, B => n623, Y => n621);
   U554 : na210 port map( A => n425, B => n624, Y => n616);
   U555 : iv110 port map( A => n501, Y => n615);
   U556 : na210 port map( A => n625, B => n544, Y => n501);
   U557 : na210 port map( A => n469, B => n481, Y => n544);
   U558 : na210 port map( A => n480, B => n472, Y => n625);
   U559 : na210 port map( A => n626, B => n627, Y => n613);
   U560 : na210 port map( A => n622, B => n586, Y => n627);
   U561 : iv110 port map( A => n628, Y => n626);
   U562 : no310 port map( A => n629, B => n630, C => n631, Y => n594);
   U563 : no210 port map( A => n620, B => n561, Y => n631);
   U564 : no210 port map( A => n534, B => n424, Y => n630);
   U565 : no210 port map( A => n487, B => n508, Y => n629);
   U566 : no310 port map( A => n632, B => n633, C => n634, Y => n593);
   U567 : no210 port map( A => n581, B => n571, Y => n634);
   U568 : no210 port map( A => n585, B => n468, Y => n633);
   U569 : na310 port map( A => n635, B => n636, C => n637, Y => rom_d(11));
   U570 : no310 port map( A => n638, B => n438, C => n614, Y => n637);
   U571 : na210 port map( A => n639, B => n640, Y => n614);
   U572 : na210 port map( A => n509, B => n641, Y => n640);
   U573 : na210 port map( A => n481, B => n562, Y => n639);
   U574 : na310 port map( A => n642, B => n643, C => n644, Y => n638);
   U575 : na210 port map( A => n469, B => n536, Y => n644);
   U576 : na210 port map( A => n645, B => n511, Y => n643);
   U577 : na210 port map( A => n624, B => n450, Y => n642);
   U578 : no210 port map( A => n552, B => n564, Y => n636);
   U579 : na210 port map( A => n646, B => n647, Y => n564);
   U580 : na210 port map( A => n623, B => n481, Y => n647);
   U581 : na210 port map( A => n612, B => n641, Y => n646);
   U582 : na210 port map( A => n648, B => n649, Y => n552);
   U583 : na210 port map( A => n449, B => n650, Y => n649);
   U584 : na210 port map( A => n457, B => n479, Y => n650);
   U585 : na210 port map( A => n469, B => n510, Y => n648);
   U586 : no210 port map( A => n651, B => n652, Y => n635);
   U587 : na310 port map( A => n653, B => n654, C => n655, Y => rom_d(10));
   U588 : iv110 port map( A => n656, Y => n655);
   U589 : na310 port map( A => n657, B => n490, C => n658, Y => n656);
   U590 : iv110 port map( A => n529, Y => n490);
   U591 : na210 port map( A => n659, B => n660, Y => n529);
   U592 : na210 port map( A => n559, B => n451, Y => n660);
   U593 : na210 port map( A => n661, B => n445, Y => n659);
   U594 : no210 port map( A => n651, B => n599, Y => n657);
   U595 : na210 port map( A => n662, B => n663, Y => n599);
   U596 : na210 port map( A => n450, B => n451, Y => n663);
   U597 : na210 port map( A => n425, B => n664, Y => n662);
   U598 : na310 port map( A => n665, B => n666, C => n667, Y => n651);
   U599 : no310 port map( A => n668, B => n669, C => n670, Y => n667);
   U600 : no210 port map( A => n482, B => n671, Y => n670);
   U601 : no210 port map( A => n672, B => n466, Y => n669);
   U602 : na310 port map( A => n673, B => n674, C => n675, Y => n668);
   U603 : na210 port map( A => n510, B => n450, Y => n675);
   U604 : na210 port map( A => n470, B => n536, Y => n674);
   U605 : na210 port map( A => n466, B => n495, Y => n470);
   U606 : na210 port map( A => n472, B => n511, Y => n673);
   U607 : no210 port map( A => n496, B => n463, Y => n666);
   U608 : no210 port map( A => n585, B => n581, Y => n463);
   U609 : no210 port map( A => n424, B => n444, Y => n496);
   U610 : no210 port map( A => n632, B => n528, Y => n665);
   U611 : na210 port map( A => n676, B => n677, Y => n528);
   U612 : na210 port map( A => n559, B => n664, Y => n677);
   U613 : na210 port map( A => n480, B => n425, Y => n676);
   U614 : no210 port map( A => n515, B => n507, Y => n632);
   U615 : no210 port map( A => n678, B => n428, Y => n654);
   U616 : na310 port map( A => n679, B => n680, C => n681, Y => n428);
   U617 : no310 port map( A => n682, B => n543, C => n600, Y => n681);
   U618 : na310 port map( A => n683, B => n684, C => n685, Y => n600);
   U619 : no210 port map( A => n686, B => n687, Y => n685);
   U620 : no210 port map( A => n688, B => n558, Y => n687);
   U621 : no310 port map( A => n623, B => n472, C => n612, Y => n688);
   U622 : no210 port map( A => n689, B => n507, Y => n686);
   U623 : no210 port map( A => n559, B => n452, Y => n689);
   U624 : na210 port map( A => n661, B => n609, Y => n684);
   U625 : iv110 port map( A => n439, Y => n683);
   U626 : na210 port map( A => n690, B => n691, Y => n439);
   U627 : na210 port map( A => n469, B => n445, Y => n691);
   U628 : na210 port map( A => n480, B => n612, Y => n690);
   U629 : na210 port map( A => n692, B => n693, Y => n543);
   U630 : na210 port map( A => n449, B => n694, Y => n693);
   U631 : na310 port map( A => n695, B => n515, C => n577, Y => n694);
   U632 : no210 port map( A => n425, B => n450, Y => n577);
   U633 : na210 port map( A => n510, B => n592, Y => n692);
   U634 : na210 port map( A => n696, B => n697, Y => n682);
   U635 : na210 port map( A => n449, B => n698, Y => n697);
   U636 : na310 port map( A => n495, B => n508, C => n576, Y => n698);
   U637 : na210 port map( A => n510, B => n699, Y => n696);
   U638 : iv110 port map( A => n700, Y => n680);
   U639 : no210 port map( A => n591, B => n438, Y => n679);
   U640 : na310 port map( A => n701, B => n702, C => n703, Y => n438);
   U641 : no210 port map( A => n704, B => n705, Y => n703);
   U642 : no210 port map( A => n456, B => n479, Y => n705);
   U643 : no210 port map( A => n483, B => n482, Y => n704);
   U644 : no210 port map( A => n425, B => n622, Y => n483);
   U645 : iv110 port map( A => n706, Y => n425);
   U646 : na210 port map( A => n641, B => n707, Y => n702);
   U647 : na210 port map( A => n585, B => n495, Y => n707);
   U648 : na210 port map( A => n451, B => n517, Y => n701);
   U649 : na210 port map( A => n515, B => n571, Y => n517);
   U650 : na210 port map( A => n708, B => n709, Y => n591);
   U651 : na210 port map( A => n586, B => n710, Y => n709);
   U652 : na210 port map( A => n479, B => n585, Y => n710);
   U653 : na210 port map( A => n471, B => n623, Y => n708);
   U654 : no210 port map( A => n437, B => n537, Y => n653);
   U655 : na210 port map( A => n711, B => n712, Y => n437);
   U656 : na210 port map( A => n586, B => n713, Y => n712);
   U657 : na310 port map( A => n714, B => n706, C => n576, Y => n713);
   U658 : iv110 port map( A => n699, Y => n576);
   U659 : na310 port map( A => n715, B => n716, C => n717, Y => rom_d(0));
   U660 : no310 port map( A => n718, B => n537, C => n652, Y => n717);
   U661 : na310 port map( A => n719, B => n720, C => n721, Y => n652);
   U662 : no310 port map( A => n722, B => n723, C => n724, Y => n721);
   U663 : no210 port map( A => n558, B => n495, Y => n724);
   U664 : no210 port map( A => n527, B => n458, Y => n723);
   U665 : na210 port map( A => n725, B => n726, Y => n722);
   U666 : na210 port map( A => n449, B => n727, Y => n726);
   U667 : na310 port map( A => n671, B => n571, C => n728, Y => n727);
   U668 : na210 port map( A => n451, B => n729, Y => n725);
   U669 : na310 port map( A => n479, B => n620, C => n495, Y => n729);
   U670 : no210 port map( A => n730, B => n731, Y => n720);
   U671 : no210 port map( A => n482, B => n714, Y => n731);
   U672 : no210 port map( A => n672, B => n444, Y => n730);
   U673 : iv110 port map( A => n609, Y => n672);
   U674 : no210 port map( A => n678, B => n598, Y => n719);
   U675 : na310 port map( A => n658, B => n418, C => n732, Y => n598);
   U676 : no310 port map( A => n733, B => n505, C => n500, Y => n732);
   U677 : no210 port map( A => n524, B => n706, Y => n500);
   U678 : no210 port map( A => n479, B => n458, Y => n505);
   U679 : no210 port map( A => n456, B => n571, Y => n733);
   U680 : iv110 port map( A => n734, Y => n418);
   U681 : na310 port map( A => n735, B => n736, C => n737, Y => n734);
   U682 : na210 port map( A => n641, B => n738, Y => n737);
   U683 : na210 port map( A => n451, B => n739, Y => n736);
   U684 : na210 port map( A => n457, B => n508, Y => n739);
   U685 : na210 port map( A => n450, B => n445, Y => n735);
   U686 : iv110 port map( A => n740, Y => n658);
   U687 : na310 port map( A => n741, B => n742, C => n743, Y => n740);
   U688 : na210 port map( A => n562, B => n641, Y => n743);
   U689 : na210 port map( A => n445, B => n592, Y => n742);
   U690 : na210 port map( A => n509, B => n664, Y => n741);
   U691 : no210 port map( A => n585, B => n507, Y => n678);
   U692 : na210 port map( A => n744, B => n745, Y => n537);
   U693 : na210 port map( A => n623, B => n451, Y => n745);
   U694 : iv110 port map( A => n524, Y => n451);
   U695 : na210 port map( A => n641, B => n452, Y => n744);
   U696 : iv110 port map( A => n466, Y => n452);
   U697 : na210 port map( A => n711, B => n502, Y => n718);
   U698 : iv110 port map( A => n746, Y => n502);
   U699 : na210 port map( A => n747, B => n588, Y => n746);
   U700 : na210 port map( A => n471, B => n562, Y => n588);
   U701 : iv110 port map( A => n507, Y => n471);
   U702 : na210 port map( A => n510, B => n535, Y => n747);
   U703 : iv110 port map( A => n558, Y => n510);
   U704 : iv110 port map( A => n748, Y => n711);
   U705 : na310 port map( A => n749, B => n750, C => n751, Y => n748);
   U706 : na210 port map( A => n535, B => n445, Y => n751);
   U707 : iv110 port map( A => n515, Y => n535);
   U708 : na210 port map( A => n480, B => n450, Y => n750);
   U709 : na210 port map( A => n469, B => n664, Y => n749);
   U710 : iv110 port map( A => n508, Y => n469);
   U711 : no210 port map( A => n493, B => n752, Y => n716);
   U712 : no210 port map( A => n554, B => n495, Y => n752);
   U713 : no210 port map( A => n586, B => n449, Y => n554);
   U714 : iv110 port map( A => n561, Y => n449);
   U715 : no210 port map( A => n468, B => n534, Y => n493);
   U716 : no210 port map( A => n753, B => n700, Y => n715);
   U717 : na310 port map( A => n754, B => n755, C => n756, Y => n700);
   U718 : no210 port map( A => n757, B => n758, Y => n756);
   U719 : iv110 port map( A => n759, Y => n758);
   U720 : no310 port map( A => n453, B => n628, C => n601, Y => n759);
   U721 : na310 port map( A => n760, B => n761, C => n762, Y => n601);
   U722 : no310 port map( A => n763, B => n764, C => n765, Y => n762);
   U723 : no210 port map( A => n479, B => n424, Y => n765);
   U724 : no210 port map( A => n515, B => n581, Y => n764);
   U725 : no210 port map( A => n458, B => n706, Y => n763);
   U726 : na210 port map( A => n562, B => n609, Y => n761);
   U727 : na210 port map( A => n456, B => n558, Y => n609);
   U728 : no210 port map( A => n766, B => n767, Y => n760);
   U729 : no210 port map( A => n488, B => n728, Y => n767);
   U730 : no210 port map( A => n553, B => n768, Y => n766);
   U731 : na310 port map( A => n769, B => n770, C => n771, Y => n628);
   U732 : no310 port map( A => n772, B => n773, C => n774, Y => n771);
   U733 : no210 port map( A => n468, B => n671, Y => n774);
   U734 : no210 port map( A => n466, B => n581, Y => n773);
   U735 : iv110 port map( A => n775, Y => n772);
   U736 : no210 port map( A => n776, B => n777, Y => n775);
   U737 : no210 port map( A => n768, B => n488, Y => n777);
   U738 : no210 port map( A => n738, B => n509, Y => n768);
   U739 : no210 port map( A => n607, B => n553, Y => n776);
   U740 : no210 port map( A => n778, B => n622, Y => n607);
   U741 : iv110 port map( A => n495, Y => n622);
   U742 : na210 port map( A => n738, B => n664, Y => n770);
   U743 : iv110 port map( A => n620, Y => n738);
   U744 : no210 port map( A => n779, B => n780, Y => n769);
   U745 : no210 port map( A => n482, B => n781, Y => n780);
   U746 : no210 port map( A => n458, B => n444, Y => n779);
   U747 : na310 port map( A => n782, B => n783, C => n784, Y => n453);
   U748 : no210 port map( A => n785, B => n786, Y => n784);
   U749 : no210 port map( A => n706, B => n558, Y => n786);
   U750 : no210 port map( A => n458, B => n457, Y => n785);
   U751 : na210 port map( A => n586, B => n645, Y => n783);
   U752 : na210 port map( A => n457, B => n571, Y => n645);
   U753 : iv110 port map( A => n468, Y => n586);
   U754 : na310 port map( A => n787, B => n788, C => rom_a(7), Y => n468);
   U755 : na210 port map( A => n612, B => n445, Y => n782);
   U756 : iv110 port map( A => n482, Y => n445);
   U757 : na310 port map( A => n789, B => n790, C => n791, Y => n757);
   U758 : na210 port map( A => n612, B => n624, Y => n791);
   U759 : iv110 port map( A => n424, Y => n624);
   U760 : iv110 port map( A => n571, Y => n612);
   U761 : na210 port map( A => n792, B => n793, Y => n571);
   U762 : na210 port map( A => n559, B => n481, Y => n790);
   U763 : iv110 port map( A => n581, Y => n481);
   U764 : iv110 port map( A => n459, Y => n559);
   U765 : na210 port map( A => n480, B => n778, Y => n789);
   U766 : iv110 port map( A => n487, Y => n480);
   U767 : no310 port map( A => n794, B => n795, C => n796, Y => n755);
   U768 : no210 port map( A => n797, B => n482, Y => n796);
   U769 : na210 port map( A => n787, B => n798, Y => n482);
   U770 : no210 port map( A => n472, B => n699, Y => n797);
   U771 : na210 port map( A => n620, B => n459, Y => n699);
   U772 : na210 port map( A => n793, B => n799, Y => n459);
   U773 : na210 port map( A => n800, B => n799, Y => n620);
   U774 : iv110 port map( A => n479, Y => n472);
   U775 : na210 port map( A => n792, B => n800, Y => n479);
   U776 : no210 port map( A => n801, B => n524, Y => n795);
   U777 : na210 port map( A => n802, B => n803, Y => n524);
   U778 : iv110 port map( A => n804, Y => n801);
   U779 : na210 port map( A => n695, B => n728, Y => n804);
   U780 : no210 port map( A => n562, B => n592, Y => n728);
   U781 : iv110 port map( A => n585, Y => n592);
   U782 : na210 port map( A => n799, B => n805, Y => n585);
   U783 : iv110 port map( A => n781, Y => n562);
   U784 : na210 port map( A => n800, B => n806, Y => n781);
   U785 : no210 port map( A => n509, B => n778, Y => n695);
   U786 : iv110 port map( A => n444, Y => n778);
   U787 : na210 port map( A => n792, B => n805, Y => n444);
   U788 : iv110 port map( A => n714, Y => n509);
   U789 : na210 port map( A => n807, B => n805, Y => n714);
   U790 : na210 port map( A => n808, B => n809, Y => n794);
   U791 : na210 port map( A => n664, B => n810, Y => n809);
   U792 : na210 port map( A => n527, B => n495, Y => n810);
   U793 : na210 port map( A => n800, B => n807, Y => n495);
   U794 : no210 port map( A => n811, B => n812, Y => n800);
   U795 : no210 port map( A => n623, B => n450, Y => n527);
   U796 : iv110 port map( A => n534, Y => n450);
   U797 : na210 port map( A => n793, B => n807, Y => n534);
   U798 : iv110 port map( A => n456, Y => n664);
   U799 : na210 port map( A => n798, B => n803, Y => n456);
   U800 : na210 port map( A => n641, B => n813, Y => n808);
   U801 : na210 port map( A => n515, B => n508, Y => n813);
   U802 : na210 port map( A => n814, B => n799, Y => n508);
   U803 : no210 port map( A => n815, B => rom_a(2), Y => n799);
   U804 : na210 port map( A => n814, B => n806, Y => n515);
   U805 : iv110 port map( A => n458, Y => n641);
   U806 : na310 port map( A => n798, B => n816, C => rom_a(6), Y => n458);
   U807 : no310 port map( A => n817, B => n818, C => n819, Y => n754);
   U808 : no210 port map( A => n553, B => n706, Y => n819);
   U809 : na210 port map( A => n792, B => n814, Y => n706);
   U810 : no210 port map( A => rom_a(3), B => rom_a(2), Y => n792);
   U811 : iv110 port map( A => n511, Y => n553);
   U812 : na210 port map( A => n581, B => n507, Y => n511);
   U813 : na310 port map( A => rom_a(5), B => n798, C => rom_a(6), Y => n507);
   U814 : no210 port map( A => n788, B => rom_a(7), Y => n798);
   U815 : na210 port map( A => n802, B => n787, Y => n581);
   U816 : no210 port map( A => n816, B => rom_a(6), Y => n787);
   U817 : no210 port map( A => n488, B => n578, Y => n818);
   U818 : no210 port map( A => n661, B => n623, Y => n578);
   U819 : iv110 port map( A => n671, Y => n623);
   U820 : na210 port map( A => n793, B => n806, Y => n671);
   U821 : no210 port map( A => rom_a(1), B => rom_a(0), Y => n793);
   U822 : iv110 port map( A => n457, Y => n661);
   U823 : iv110 port map( A => n536, Y => n488);
   U824 : na210 port map( A => n487, B => n424, Y => n536);
   U825 : na310 port map( A => n802, B => n816, C => rom_a(6), Y => n424);
   U826 : iv110 port map( A => rom_a(5), Y => n816);
   U827 : na310 port map( A => n802, B => rom_a(5), C => rom_a(6), Y => n487);
   U828 : no210 port map( A => rom_a(7), B => rom_a(4), Y => n802);
   U829 : no210 port map( A => n466, B => n561, Y => n817);
   U830 : na310 port map( A => n803, B => rom_a(4), C => rom_a(7), Y => n561);
   U831 : na210 port map( A => n806, B => n805, Y => n466);
   U832 : no210 port map( A => n812, B => rom_a(1), Y => n805);
   U833 : iv110 port map( A => rom_a(0), Y => n812);
   U834 : no210 port map( A => n820, B => n815, Y => n806);
   U835 : iv110 port map( A => rom_a(3), Y => n815);
   U836 : no210 port map( A => n457, B => n558, Y => n753);
   U837 : na310 port map( A => n803, B => n788, C => rom_a(7), Y => n558);
   U838 : iv110 port map( A => rom_a(4), Y => n788);
   U839 : no210 port map( A => rom_a(6), B => rom_a(5), Y => n803);
   U840 : na210 port map( A => n807, B => n814, Y => n457);
   U841 : no210 port map( A => n811, B => rom_a(0), Y => n814);
   U842 : iv110 port map( A => rom_a(1), Y => n811);
   U843 : no210 port map( A => n820, B => rom_a(3), Y => n807);
   U844 : iv110 port map( A => rom_a(2), Y => n820);

end synthesised;



