configuration reg_o_behaviour_cfg of reg_o is
   for behaviour
   end for;
end reg_o_behaviour_cfg;


