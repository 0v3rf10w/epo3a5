configuration reg_6_behaviour_cfg of reg_6 is
   for behaviour
   end for;
end reg_6_behaviour_cfg;


