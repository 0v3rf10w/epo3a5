configuration stream_behaviour_cfg of stream is
   for behaviour
   end for;
end stream_behaviour_cfg;


