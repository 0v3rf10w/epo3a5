configuration buf_arg_behaviour_cfg of buf_arg is
   for behaviour
   end for;
end buf_arg_behaviour_cfg;


