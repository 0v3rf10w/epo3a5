library IEEE;
use IEEE.std_logic_1164.all;

entity ROM is
port
(
    rom_a:    in std_logic_vector (7 DOWNTO 0);     -- address
    rom_d:    out std_logic_vector (11 DOWNTO 0)    -- instruction
);
end ROM;

architecture behavioural OF ROM IS
begin
    with rom_a select
    rom_d <=
"111100000000" when "00000000",
"011000000001" when "00000001",
"101000101111" when "00000010",
"100000000001" when "00000011",
"010000001110" when "00000100",
"011000000001" when "00000101",
"101000011111" when "00000110",
"100000000001" when "00000111",
"010000110010" when "00001000",
"011000000001" when "00001001",
"101000001111" when "00001010",
"100000000001" when "00001011",
"010001011001" when "00001100",
"000100000000" when "00001101",
"111100000000" when "00001110",
"011000000001" when "00001111",
"101000101111" when "00010000",
"100000000001" when "00010001",
"010000001110" when "00010010",
"111100000000" when "00010011",
"011000000001" when "00010100",
"110000001111" when "00010101",
"011100000010" when "00010110",
"011000000001" when "00010111",
"110000010000" when "00011000",
"001100011100" when "00011001",
"010100000001" when "00011010",
"011100000011" when "00011011",
"011000000001" when "00011100",
"110000100000" when "00011101",
"001100100010" when "00011110",
"011000000011" when "00011111",
"100000000010" when "00100000",
"011100000011" when "00100001",
"011000000001" when "00100010",
"110001000000" when "00100011",
"001100101000" when "00100100",
"011000000011" when "00100101",
"100000000100" when "00100110",
"011100000011" when "00100111",
"011000000001" when "00101000",
"110010000000" when "00101001",
"001100101110" when "00101010",
"011000000011" when "00101011",
"100000001000" when "00101100",
"011100000011" when "00101101",
"011000000011" when "00101110",
"100100000010" when "00101111",
"011100000001" when "00110000",
"000100000000" when "00110001",
"111100000000" when "00110010",
"011000000001" when "00110011",
"101000011111" when "00110100",
"100000000001" when "00110101",
"010000110010" when "00110110",
"111100000000" when "00110111",
"011000000001" when "00111000",
"110000001111" when "00111001",
"011100000010" when "00111010",
"011000000001" when "00111011",
"110000010000" when "00111100",
"001101000000" when "00111101",
"010100000001" when "00111110",
"011100000011" when "00111111",
"011000000001" when "01000000",
"110000100000" when "01000001",
"001101000110" when "01000010",
"011000000011" when "01000011",
"100000000010" when "01000100",
"011100000011" when "01000101",
"011000000001" when "01000110",
"110001000000" when "01000111",
"001101001100" when "01001000",
"011000000011" when "01001001",
"100000000100" when "01001010",
"011100000011" when "01001011",
"011000000001" when "01001100",
"110010000000" when "01001101",
"001101010010" when "01001110",
"011000000011" when "01001111",
"100000001000" when "01010000",
"011100000011" when "01010001",
"011000000011" when "01010010",
"101011111111" when "01010011",
"100000000001" when "01010100",
"100100000010" when "01010101",
"011100000001" when "01010110",
"111100000000" when "01010111",
"000100000000" when "01011000",
"111100000000" when "01011001",
"011000000001" when "01011010",
"101000001111" when "01011011",
"100000000001" when "01011100",
"010001011001" when "01011101",
"011000000001" when "01011110",
"110000001111" when "01011111",
"011100000010" when "01100000",
"011000000001" when "01100001",
"110000010000" when "01100010",
"001101100110" when "01100011",
"010100000001" when "01100100",
"011100000011" when "01100101",
"011000000001" when "01100110",
"110000100000" when "01100111",
"001101101100" when "01101000",
"011000000011" when "01101001",
"100000000010" when "01101010",
"011100000011" when "01101011",
"011000000001" when "01101100",
"110001000000" when "01101101",
"001101110010" when "01101110",
"011000000011" when "01101111",
"100000000100" when "01110000",
"011100000011" when "01110001",
"011000000001" when "01110010",
"110010000000" when "01110011",
"001101111000" when "01110100",
"011000000011" when "01110101",
"100000001000" when "01110110",
"011100000011" when "01110111",
"011000000010" when "01111000",
"110000000001" when "01111001",
"001110100010" when "01111010",
"011000000011" when "01111011",
"011100000100" when "01111100",
"011000000010" when "01111101",
"110000000010" when "01111110",
"001110100101" when "01111111",
"011000000010" when "10000000",
"100100000011" when "10000001",
"011100000101" when "10000010",
"011000000010" when "10000011",
"110000000100" when "10000100",
"001110101000" when "10000101",
"011000000011" when "10000110",
"100100000011" when "10000111",
"011100001000" when "10001000",
"011000001000" when "10001001",
"100100001000" when "10001010",
"011100000110" when "10001011",
"011000000010" when "10001100",
"110000001000" when "10001101",
"001110101011" when "10001110",
"011000000011" when "10001111",
"100100000011" when "10010000",
"011100001000" when "10010001",
"011000001000" when "10010010",
"100100001000" when "10010011",
"011100001000" when "10010100",
"011000001000" when "10010101",
"100100001000" when "10010110",
"011100000111" when "10010111",
"011000000100" when "10011000",
"100100000101" when "10011001",
"011100001000" when "10011010",
"011000000110" when "10011011",
"100100000111" when "10011100",
"011100001001" when "10011101",
"011000001000" when "10011110",
"100100001001" when "10011111",
"011100000001" when "10100000",
"000100000000" when "10100001",
"010100000000" when "10100010",
"011100000100" when "10100011",
"000101111101" when "10100100",
"010100000000" when "10100101",
"011100000101" when "10100110",
"000110000011" when "10100111",
"010100000000" when "10101000",
"011100000110" when "10101001",
"000110001100" when "10101010",
"010100000000" when "10101011",
"011100000111" when "10101100",
"000110011000" when "10101101",



"000000000000" when others;
end behavioural;

