configuration vidcounter_behavioural_cfg of vidcounter is
   for behavioural
   end for;
end vidcounter_behavioural_cfg;


