configuration reg_7_behaviour_cfg of reg_7 is
   for behaviour
   end for;
end reg_7_behaviour_cfg;


