configuration blackbox_synthesised_cfg of blackbox is
   for synthesised
      for all: stream use configuration work.stream_behaviour_cfg;
      end for;
   end for;
end blackbox_synthesised_cfg;


