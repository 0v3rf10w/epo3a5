library IEEE;
use IEEE.std_logic_1164.ALL;

entity tbuf40_tb is
end tbuf40_tb;


