configuration tbuf_tb_behaviour_cfg of tbuf_tb is
   for behaviour
      for all: tbuf use configuration work.tbuf_behaviour_cfg;
      end for;
   end for;
end tbuf_tb_behaviour_cfg;


