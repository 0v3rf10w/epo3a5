configuration spi_extracted_cfg of spi is
   for extracted
   end for;
end spi_extracted_cfg;


