configuration sdcard_behavioural_cfg of sdcard is
   for behavioural
   end for;
end sdcard_behavioural_cfg;


