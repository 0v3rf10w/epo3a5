configuration klokdeler_extracted_cfg of klokdeler is
   for extracted
   end for;
end klokdeler_extracted_cfg;


