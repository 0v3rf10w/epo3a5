configuration dff_behavioural_cfg of dff is
   for behavioural
   end for;
end dff_behavioural_cfg;


