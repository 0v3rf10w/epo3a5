library IEEE;
use IEEE.std_logic_1164.ALL;

entity tbuf is
   port(A :in    std_logic;
        Y:out   std_logic;
        E      :in    std_logic);
end tbuf;


