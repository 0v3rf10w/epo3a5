library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of iv is
begin
Y <= not A;
end behaviour;


