configuration stream_behaviour_cfg of stream is
   for behaviour
      for all: tbuf use configuration work.tbuf_behaviour_cfg;
      end for;
   end for;
end stream_behaviour_cfg;


