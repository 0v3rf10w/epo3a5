configuration buf_i_behaviour_cfg of buf_i is
   for behaviour
   end for;
end buf_i_behaviour_cfg;


