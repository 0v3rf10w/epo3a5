configuration reg_cluster_behavioural_cfg of reg_cluster is
   for behavioural
      for all: reg_o use configuration work.reg_o_behaviour_cfg;
      end for;
      for all: reg_2 use configuration work.reg_2_behaviour_cfg;
      end for;
      for all: reg_3 use configuration work.reg_3_behaviour_cfg;
      end for;
      for all: reg_4 use configuration work.reg_4_behaviour_cfg;
      end for;
      for all: reg_5 use configuration work.reg_5_behaviour_cfg;
      end for;
      for all: reg_6 use configuration work.reg_6_behaviour_cfg;
      end for;
      for all: reg_7 use configuration work.reg_7_behaviour_cfg;
      end for;
      for all: reg_8 use configuration work.reg_8_behaviour_cfg;
      end for;
      for all: reg_9 use configuration work.reg_9_behaviour_cfg;
      end for;
      for all: reg_10 use configuration work.reg_10_behaviour_cfg;
      end for;
      for all: buf_i use configuration work.buf_i_behaviour_cfg;
      end for;
      for all: buf_2 use configuration work.buf_2_behaviour_cfg;
      end for;
      for all: buf_3 use configuration work.buf_3_behaviour_cfg;
      end for;
      for all: buf_4 use configuration work.buf_4_behaviour_cfg;
      end for;
      for all: buf_5 use configuration work.buf_5_behaviour_cfg;
      end for;
      for all: buf_6 use configuration work.buf_6_behaviour_cfg;
      end for;
      for all: buf_7 use configuration work.buf_7_behaviour_cfg;
      end for;
      for all: buf_8 use configuration work.buf_8_behaviour_cfg;
      end for;
      for all: buf_9 use configuration work.buf_9_behaviour_cfg;
      end for;
      for all: buf_10 use configuration work.buf_10_behaviour_cfg;
      end for;
   end for;
end reg_cluster_behavioural_cfg;


