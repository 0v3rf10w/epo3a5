configuration spi_tb_structural_cfg of spi_tb is
   for structural
      for all: spi use configuration work.spi_structural_cfg;
      end for;
   end for;
end spi_tb_structural_cfg;


