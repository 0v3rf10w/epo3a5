configuration blackbox_extracted_cfg of blackbox is
   for extracted
   end for;
end blackbox_extracted_cfg;


