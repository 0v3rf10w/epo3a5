library IEEE;
use IEEE.std_logic_1164.ALL;

entity dff is
   port(clk :in    std_logic;
        d   :in    std_logic;
reset : in std_logic;
        q   :out   std_logic;
        qbar:out   std_logic);
end dff;









