configuration buf_10_behaviour_cfg of buf_10 is
   for behaviour
   end for;
end buf_10_behaviour_cfg;


