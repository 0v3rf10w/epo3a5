configuration buf_2_behaviour_cfg of buf_2 is
   for behaviour
   end for;
end buf_2_behaviour_cfg;


