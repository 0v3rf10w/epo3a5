configuration reg_a_behaviour_cfg of reg_a is
   for behaviour
   end for;
end reg_a_behaviour_cfg;


