configuration tbuf_behaviour_cfg of tbuf is
   for behaviour
   end for;
end tbuf_behaviour_cfg;


