configuration pc_counter_behaviour_cfg of pc_counter is
   for behaviour
   end for;
end pc_counter_behaviour_cfg;


