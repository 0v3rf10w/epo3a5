configuration tbdff_behavioural_cfg of tbdff is
   for behavioural
      for all: dff use configuration work.dff_behavioural_cfg;
      end for;
   end for;
end tbdff_behavioural_cfg;


