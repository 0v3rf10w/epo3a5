configuration reg_8_behaviour_cfg of reg_8 is
   for behaviour
   end for;
end reg_8_behaviour_cfg;


