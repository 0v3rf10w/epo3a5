configuration iv_behaviour_cfg of iv is
   for behaviour
   end for;
end iv_behaviour_cfg;


