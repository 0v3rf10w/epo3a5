library IEEE;
use IEEE.std_logic_1164.ALL;

entity stream_tb is
end stream_tb;


