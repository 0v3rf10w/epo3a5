configuration control_behavioural_cfg of control is
   for behavioural
   end for;
end control_behavioural_cfg;


