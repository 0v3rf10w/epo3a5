configuration buf_4_behaviour_cfg of buf_4 is
   for behaviour
   end for;
end buf_4_behaviour_cfg;


