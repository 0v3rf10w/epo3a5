configuration buf_a_behaviour_cfg of buf_a is
   for behaviour
   end for;
end buf_a_behaviour_cfg;


