configuration gate_behavioral_cfg of gate is
   for behavioral
   end for;
end gate_behavioral_cfg;


