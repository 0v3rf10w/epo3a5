configuration shift_reg_behavioral_cfg of shift_reg is
   for behavioral
   end for;
end shift_reg_behavioral_cfg;


