configuration shift_reg_structural_cfg of shift_reg is
   for structural
   end for;
end shift_reg_structural_cfg;


