configuration vsync_behaviour_cfg of vsync is
   for behaviour
   end for;
end vsync_behaviour_cfg;


