configuration instr_buf_behaviour_cfg of instr_buf is
   for behaviour
   end for;
end instr_buf_behaviour_cfg;


