configuration stream_tb_behaviour_cfg of stream_tb is
   for behaviour
      for all: stream use configuration work.stream_behaviour_cfg;
      end for;
   end for;
end stream_tb_behaviour_cfg;


