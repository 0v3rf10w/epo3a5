configuration tb_behaviouralexta_cfg of tb is
   for behavioural
      for all: klokdeler use configuration work.klokdeler_extracted_cfg;
      end for;
   end for;
end tb_behaviouralexta_cfg;


