configuration buf_8_behaviour_cfg of buf_8 is
   for behaviour
   end for;
end buf_8_behaviour_cfg;


